-- Testbench automatically generated online
-- at https://vhdl.lapinoo.net
-- Generation date : 15.10.2020 13:05:38 UTC

library ieee;
use ieee.std_logic_1164.all;

entity tb_and_gate is
end tb_and_gate;

architecture tb of tb_and_gate is

    component and_gate
        port (a : in std_logic;
              b : in std_logic;
              c : out std_logic);
    end component;

    signal a : std_logic;
    signal b : std_logic;
    signal c : std_logic;

begin

    dut : and_gate
    port map (a => a,
              b => b,
              c => c);

    stimuli : process
    begin
        -- EDIT Adapt initialization as needed
        a <= '0';
        b <= '0';
        wait for 10 ns;
        
        a <= '0';
        b <= '1';
        wait for 10 ns;
        
        a <= '1';
        b <= '1'; 
        
        wait;
    end process;

end tb;


